library verilog;
use verilog.vl_types.all;
entity ddr2_phy_init is
    generic(
        BANK_WIDTH      : integer := 2;
        CKE_WIDTH       : integer := 1;
        COL_WIDTH       : integer := 10;
        CS_BITS         : integer := 0;
        CS_NUM          : integer := 1;
        DQ_WIDTH        : integer := 72;
        ODT_WIDTH       : integer := 1;
        ROW_WIDTH       : integer := 14;
        ADDITIVE_LAT    : integer := 0;
        BURST_LEN       : integer := 4;
        TWO_T_TIME_EN   : integer := 0;
        BURST_TYPE      : integer := 0;
        CAS_LAT         : integer := 5;
        ODT_TYPE        : integer := 1;
        REDUCE_DRV      : integer := 0;
        REG_ENABLE      : integer := 1;
        TWR             : integer := 15000;
        CLK_PERIOD      : integer := 3000;
        DDR_TYPE        : integer := 1;
        SIM_ONLY        : integer := 0
    );
    port(
        clk0            : in     vl_logic;
        clkdiv0         : in     vl_logic;
        rst0            : in     vl_logic;
        rstdiv0         : in     vl_logic;
        calib_done      : in     vl_logic_vector(3 downto 0);
        ctrl_ref_flag   : in     vl_logic;
        calib_ref_req   : in     vl_logic;
        calib_start     : out    vl_logic_vector(3 downto 0);
        calib_ref_done  : out    vl_logic;
        phy_init_wren   : out    vl_logic;
        phy_init_rden   : out    vl_logic;
        phy_init_addr   : out    vl_logic_vector;
        phy_init_ba     : out    vl_logic_vector;
        phy_init_ras_n  : out    vl_logic;
        phy_init_cas_n  : out    vl_logic;
        phy_init_we_n   : out    vl_logic;
        phy_init_cs_n   : out    vl_logic_vector;
        phy_init_cke    : out    vl_logic_vector;
        phy_init_done   : out    vl_logic;
        phy_init_data_sel: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CKE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CS_BITS : constant is 1;
    attribute mti_svvh_generic_type of CS_NUM : constant is 1;
    attribute mti_svvh_generic_type of DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ADDITIVE_LAT : constant is 1;
    attribute mti_svvh_generic_type of BURST_LEN : constant is 1;
    attribute mti_svvh_generic_type of TWO_T_TIME_EN : constant is 1;
    attribute mti_svvh_generic_type of BURST_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CAS_LAT : constant is 1;
    attribute mti_svvh_generic_type of ODT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of REDUCE_DRV : constant is 1;
    attribute mti_svvh_generic_type of REG_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TWR : constant is 1;
    attribute mti_svvh_generic_type of CLK_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of DDR_TYPE : constant is 1;
    attribute mti_svvh_generic_type of SIM_ONLY : constant is 1;
end ddr2_phy_init;
