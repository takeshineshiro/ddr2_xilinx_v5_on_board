library verilog;
use verilog.vl_types.all;
entity ddr2_phy_calib is
    generic(
        DQ_WIDTH        : integer := 72;
        DQ_BITS         : integer := 7;
        DQ_PER_DQS      : integer := 8;
        DQS_BITS        : integer := 4;
        DQS_WIDTH       : integer := 9;
        ADDITIVE_LAT    : integer := 0;
        CAS_LAT         : integer := 5;
        REG_ENABLE      : integer := 1;
        CLK_PERIOD      : integer := 3000;
        SIM_ONLY        : integer := 0;
        DEBUG_EN        : integer := 0
    );
    port(
        clk             : in     vl_logic;
        clkdiv          : in     vl_logic;
        rstdiv          : in     vl_logic;
        calib_start     : in     vl_logic_vector(3 downto 0);
        ctrl_rden       : in     vl_logic;
        phy_init_rden   : in     vl_logic;
        rd_data_rise    : in     vl_logic_vector;
        rd_data_fall    : in     vl_logic_vector;
        calib_ref_done  : in     vl_logic;
        calib_done      : out    vl_logic_vector(3 downto 0);
        calib_ref_req   : out    vl_logic;
        calib_rden      : out    vl_logic_vector;
        calib_rden_sel  : out    vl_logic_vector;
        dlyrst_dq       : out    vl_logic;
        dlyce_dq        : out    vl_logic_vector;
        dlyinc_dq       : out    vl_logic_vector;
        dlyrst_dqs      : out    vl_logic;
        dlyce_dqs       : out    vl_logic_vector;
        dlyinc_dqs      : out    vl_logic_vector;
        dlyrst_gate     : out    vl_logic_vector;
        dlyce_gate      : out    vl_logic_vector;
        dlyinc_gate     : out    vl_logic_vector;
        en_dqs          : out    vl_logic_vector;
        rd_data_sel     : out    vl_logic_vector;
        dbg_idel_up_all : in     vl_logic;
        dbg_idel_down_all: in     vl_logic;
        dbg_idel_up_dq  : in     vl_logic;
        dbg_idel_down_dq: in     vl_logic;
        dbg_idel_up_dqs : in     vl_logic;
        dbg_idel_down_dqs: in     vl_logic;
        dbg_idel_up_gate: in     vl_logic;
        dbg_idel_down_gate: in     vl_logic;
        dbg_sel_idel_dq : in     vl_logic_vector;
        dbg_sel_all_idel_dq: in     vl_logic;
        dbg_sel_idel_dqs: in     vl_logic_vector;
        dbg_sel_all_idel_dqs: in     vl_logic;
        dbg_sel_idel_gate: in     vl_logic_vector;
        dbg_sel_all_idel_gate: in     vl_logic;
        dbg_calib_done  : out    vl_logic_vector(3 downto 0);
        dbg_calib_err   : out    vl_logic_vector(3 downto 0);
        dbg_calib_dq_tap_cnt: out    vl_logic_vector;
        dbg_calib_dqs_tap_cnt: out    vl_logic_vector;
        dbg_calib_gate_tap_cnt: out    vl_logic_vector;
        dbg_calib_rd_data_sel: out    vl_logic_vector;
        dbg_calib_rden_dly: out    vl_logic_vector;
        dbg_calib_gate_dly: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DQ_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQ_PER_DQS : constant is 1;
    attribute mti_svvh_generic_type of DQS_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ADDITIVE_LAT : constant is 1;
    attribute mti_svvh_generic_type of CAS_LAT : constant is 1;
    attribute mti_svvh_generic_type of REG_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CLK_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of SIM_ONLY : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_EN : constant is 1;
end ddr2_phy_calib;
